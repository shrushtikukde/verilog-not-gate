module not_gate(y,a);
  input a;
  output y;
  assign y= ~a;
endmodule
